module Instruction_Memory#(
    parameter 
)